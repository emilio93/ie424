`timescale 1ns / 1ps
module TestBench_VGAAdapter;

	// Inputs
	reg Clock;
	reg Reset;

endmodule
